`timescale 1ns / 1ps
module mackey_glass_block_16bit
(
    input [32 - 1 : 0] din,
    output reg [32 - 1 : 0] dout
);

always @(din) 
begin
    if (din <= 16'h0000) dout <= 32'h0000_0008;
    else if (din <= 16'h016C) dout <= 32'h0000_0014;
    else if (din <= 16'h02D8) dout <= 32'h0000_0046;
    else if (din <= 16'h0444) dout <= 32'h0000_0073;
    else if (din <= 16'h05B0) dout <= 32'h0000_0093;
    else if (din <= 16'h071C) dout <= 32'h0000_00C1;
    else if (din <= 16'h0888) dout <= 32'h0000_00EE;
    else if (din <= 16'h09F4) dout <= 32'h0000_010E;
    else if (din <= 16'h0B60) dout <= 32'h0000_013B;
    else if (din <= 16'h0CCC) dout <= 32'h0000_016D;
    else if (din <= 16'h0E38) dout <= 32'h0000_0189;
    else if (din <= 16'h0FA4) dout <= 32'h0000_01BA;
    else if (din <= 16'h1111) dout <= 32'h0000_01DF;
    else if (din <= 16'h127D) dout <= 32'h0000_0208;
    else if (din <= 16'h13E9) dout <= 32'h0000_0235;
    else if (din <= 16'h1555) dout <= 32'h0000_0256;
    else if (din <= 16'h16C1) dout <= 32'h0000_0283;
    else if (din <= 16'h182D) dout <= 32'h0000_02B0;
    else if (din <= 16'h1999) dout <= 32'h0000_02D1;
    else if (din <= 16'h1B05) dout <= 32'h0000_02FE;
    else if (din <= 16'h1C71) dout <= 32'h0000_032F;
    else if (din <= 16'h1DDD) dout <= 32'h0000_034C;
    else if (din <= 16'h1F49) dout <= 32'h0000_037D;
    else if (din <= 16'h20B6) dout <= 32'h0000_03AA;
    else if (din <= 16'h2222) dout <= 32'h0000_03C7;
    else if (din <= 16'h238E) dout <= 32'h0000_03F8;
    else if (din <= 16'h24FA) dout <= 32'h0000_0414;
    else if (din <= 16'h2666) dout <= 32'h0000_0446;
    else if (din <= 16'h27D2) dout <= 32'h0000_0473;
    else if (din <= 16'h293E) dout <= 32'h0000_0493;
    else if (din <= 16'h2AAA) dout <= 32'h0000_04C1;
    else if (din <= 16'h2C16) dout <= 32'h0000_04EE;
    else if (din <= 16'h2D82) dout <= 32'h0000_0537;
    else if (din <= 16'h2EEE) dout <= 32'h0000_053B;
    else if (din <= 16'h305B) dout <= 32'h0000_0568;
    else if (din <= 16'h31C7) dout <= 32'h0000_0589;
    else if (din <= 16'h3333) dout <= 32'h0000_05BA;
    else if (din <= 16'h349F) dout <= 32'h0000_05D7;
    else if (din <= 16'h360B) dout <= 32'h0000_0608;
    else if (din <= 16'h3777) dout <= 32'h0000_0635;
    else if (din <= 16'h38E3) dout <= 32'h0000_0656;
    else if (din <= 16'h3A4F) dout <= 32'h0000_0683;
    else if (din <= 16'h3BBB) dout <= 32'h0000_06B0;
    else if (din <= 16'h3D27) dout <= 32'h0000_06D1;
    else if (din <= 16'h3E93) dout <= 32'h0000_06FE;
    else if (din <= 16'h4000) dout <= 32'h0000_072B;
    else if (din <= 16'h416C) dout <= 32'h0000_074C;
    else if (din <= 16'h42D8) dout <= 32'h0000_0779;
    else if (din <= 16'h4444) dout <= 32'h0000_079A;
    else if (din <= 16'h45B0) dout <= 32'h0000_07C7;
    else if (din <= 16'h471C) dout <= 32'h0000_07F4;
    else if (din <= 16'h4888) dout <= 32'h0000_0814;
    else if (din <= 16'h49F4) dout <= 32'h0000_0842;
    else if (din <= 16'h4B60) dout <= 32'h0000_086F;
    else if (din <= 16'h4CCC) dout <= 32'h0000_088F;
    else if (din <= 16'h4E38) dout <= 32'h0000_08BC;
    else if (din <= 16'h4FA4) dout <= 32'h0000_08E9;
    else if (din <= 16'h5111) dout <= 32'h0000_090A;
    else if (din <= 16'h527D) dout <= 32'h0000_0937;
    else if (din <= 16'h53E9) dout <= 32'h0000_0954;
    else if (din <= 16'h5555) dout <= 32'h0000_0981;
    else if (din <= 16'h56C1) dout <= 32'h0000_09AE;
    else if (din <= 16'h582D) dout <= 32'h0000_09CB;
    else if (din <= 16'h5999) dout <= 32'h0000_09F8;
    else if (din <= 16'h5B05) dout <= 32'h0000_0A21;
    else if (din <= 16'h5C71) dout <= 32'h0000_0A42;
    else if (din <= 16'h5DDD) dout <= 32'h0000_0A6A;
    else if (din <= 16'h5F49) dout <= 32'h0000_0A93;
    else if (din <= 16'h60B6) dout <= 32'h0000_0AB0;
    else if (din <= 16'h6222) dout <= 32'h0000_0AD9;
    else if (din <= 16'h638E) dout <= 32'h0000_0AF2;
    else if (din <= 16'h64FA) dout <= 32'h0000_0B17;
    else if (din <= 16'h6666) dout <= 32'h0000_0B3B;
    else if (din <= 16'h67D2) dout <= 32'h0000_0B54;
    else if (din <= 16'h693E) dout <= 32'h0000_0B75;
    else if (din <= 16'h6AAA) dout <= 32'h0000_0B91;
    else if (din <= 16'h6C16) dout <= 32'h0000_0BA6;
    else if (din <= 16'h6D82) dout <= 32'h0000_0BBE;
    else if (din <= 16'h6EEE) dout <= 32'h0000_0BD7;
    else if (din <= 16'h705B) dout <= 32'h0000_0BE3;
    else if (din <= 16'h71C7) dout <= 32'h0000_0BF0;
    else if (din <= 16'h7333) dout <= 32'h0000_0BF8;
    else if (din <= 16'h749F) dout <= 32'h0000_0C00;
    else if (din <= 16'h760B) dout <= 32'h0000_0C00;
    else if (din <= 16'h7777) dout <= 32'h0000_0C00;
    else if (din <= 16'h78E3) dout <= 32'h0000_0BF4;
    else if (din <= 16'h7A4F) dout <= 32'h0000_0BE3;
    else if (din <= 16'h7BBB) dout <= 32'h0000_0BD3;
    else if (din <= 16'h7D27) dout <= 32'h0000_0BBA;
    else if (din <= 16'h7E93) dout <= 32'h0000_0B96;
    else if (din <= 16'h8000) dout <= 32'h0000_0B7D;
    else if (din <= 16'h816C) dout <= 32'h0000_0B4C;
    else if (din <= 16'h82D8) dout <= 32'h0000_0B2B;
    else if (din <= 16'h8444) dout <= 32'h0000_0AEE;
    else if (din <= 16'h85B0) dout <= 32'h0000_0AAC;
    else if (din <= 16'h871C) dout <= 32'h0000_0A7B;
    else if (din <= 16'h8888) dout <= 32'h0000_0A31;
    else if (din <= 16'h89F4) dout <= 32'h0000_09DF;
    else if (din <= 16'h8B60) dout <= 32'h0000_09A2;
    else if (din <= 16'h8CCC) dout <= 32'h0000_0948;
    else if (din <= 16'h8E38) dout <= 32'h0000_08E5;
    else if (din <= 16'h8FA4) dout <= 32'h0000_08A0;
    else if (din <= 16'h9111) dout <= 32'h0000_0835;
    else if (din <= 16'h927D) dout <= 32'h0000_07C3;
    else if (din <= 16'h93E9) dout <= 32'h0000_0775;
    else if (din <= 16'h9555) dout <= 32'h0000_06FE;
    else if (din <= 16'h96C1) dout <= 32'h0000_06A8;
    else if (din <= 16'h982D) dout <= 32'h0000_0629;
    else if (din <= 16'h9999) dout <= 32'h0000_05A2;
    else if (din <= 16'h9B05) dout <= 32'h0000_0548;
    else if (din <= 16'h9C71) dout <= 32'h0000_04BC;
    else if (din <= 16'h9DDD) dout <= 32'h0000_042D;
    else if (din <= 16'h9F49) dout <= 32'h0000_03CB;
    else if (din <= 16'hA0B6) dout <= 32'h0000_033F;
    else if (din <= 16'hA222) dout <= 32'h0000_02BC;
    else if (din <= 16'hA38E) dout <= 32'h0000_0273;
    else if (din <= 16'hA4FA) dout <= 32'h0000_021D;
    else if (din <= 16'hA666) dout <= 32'h0000_01F0;
    else if (din <= 16'hA7D2) dout <= 32'h0000_01B6;
    else if (din <= 16'hA93E) dout <= 32'h0000_0191;
    else if (din <= 16'hAAAA) dout <= 32'h0000_0175;
    else if (din <= 16'hAC16) dout <= 32'h0000_0158;
    else if (din <= 16'hAD82) dout <= 32'h0000_013F;
    else if (din <= 16'hAEEE) dout <= 32'h0000_012B;
    else if (din <= 16'hB05B) dout <= 32'h0000_011F;
    else if (din <= 16'hB1C7) dout <= 32'h0000_010A;
    else if (din <= 16'hB333) dout <= 32'h0000_0102;
    else if (din <= 16'hB49F) dout <= 32'h0000_00F6;
    else if (din <= 16'hB60B) dout <= 32'h0000_00EE;
    else if (din <= 16'hB777) dout <= 32'h0000_00E1;
    else if (din <= 16'hB8E3) dout <= 32'h0000_00D9;
    else if (din <= 16'hBA4F) dout <= 32'h0000_00CD;
    else if (din <= 16'hBBBB) dout <= 32'h0000_00C9;
    else if (din <= 16'hBD27) dout <= 32'h0000_00C1;
    else if (din <= 16'hBE93) dout <= 32'h0000_00BC;
    else if (din <= 16'hC000) dout <= 32'h0000_00B4;
    else if (din <= 16'hC16C) dout <= 32'h0000_00B0;
    else if (din <= 16'hC2D8) dout <= 32'h0000_00AC;
    else if (din <= 16'hC444) dout <= 32'h0000_00A4;
    else if (din <= 16'hC5B0) dout <= 32'h0000_00A0;
    else if (din <= 16'hC71C) dout <= 32'h0000_009C;
    else if (din <= 16'hC888) dout <= 32'h0000_0098;
    else if (din <= 16'hC9F4) dout <= 32'h0000_0093;
    else if (din <= 16'hCB60) dout <= 32'h0000_0093;
    else if (din <= 16'hCCCC) dout <= 32'h0000_008B;
    else if (din <= 16'hCE38) dout <= 32'h0000_008B;
    else if (din <= 16'hCFA4) dout <= 32'h0000_0087;
    else if (din <= 16'hD111) dout <= 32'h0000_0083;
    else if (din <= 16'hD27D) dout <= 32'h0000_0083;
    else if (din <= 16'hD3E9) dout <= 32'h0000_007F;
    else if (din <= 16'hD555) dout <= 32'h0000_007B;
    else if (din <= 16'hD6C1) dout <= 32'h0000_007B;
    else if (din <= 16'hD82D) dout <= 32'h0000_0077;
    else if (din <= 16'hD999) dout <= 32'h0000_0077;
    else if (din <= 16'hDB05) dout <= 32'h0000_0073;
    else if (din <= 16'hDC71) dout <= 32'h0000_006F;
    else if (din <= 16'hDDDD) dout <= 32'h0000_006F;
    else if (din <= 16'hDF49) dout <= 32'h0000_006A;
    else if (din <= 16'hE0B6) dout <= 32'h0000_006A;
    else if (din <= 16'hE222) dout <= 32'h0000_006A;
    else if (din <= 16'hE38E) dout <= 32'h0000_0066;
    else if (din <= 16'hE4FA) dout <= 32'h0000_0062;
    else if (din <= 16'hE666) dout <= 32'h0000_0062;
    else if (din <= 16'hE7D2) dout <= 32'h0000_0062;
    else if (din <= 16'hE93E) dout <= 32'h0000_0062;
    else if (din <= 16'hEAAA) dout <= 32'h0000_005E;
    else if (din <= 16'hEC16) dout <= 32'h0000_005E;
    else if (din <= 16'hED82) dout <= 32'h0000_005E;
    else if (din <= 16'hEEEE) dout <= 32'h0000_005A;
    else if (din <= 16'hF05B) dout <= 32'h0000_005A;
    else if (din <= 16'hF1C7) dout <= 32'h0000_005A;
    else if (din <= 16'hF333) dout <= 32'h0000_0056;
    else if (din <= 16'hF49F) dout <= 32'h0000_0056;
    else if (din <= 16'hF60B) dout <= 32'h0000_0056;
    else if (din <= 16'hF777) dout <= 32'h0000_0056;
    else if (din <= 16'hF8E3) dout <= 32'h0000_0052;
    else if (din <= 16'hFA4F) dout <= 32'h0000_0052;
    else if (din <= 16'hFBBB) dout <= 32'h0000_0052;
    else if (din <= 16'hFD27) dout <= 32'h0000_0052;
    else if (din <= 16'hFE93) dout <= 32'h0000_004E;
    else if (din <= 16'hFFFF) dout <= 32'h0000_004E;
    else dout <= 32'h0000_0000;
end


endmodule