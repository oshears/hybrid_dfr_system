`timescale 1ns / 1ps
module mackey_glass_block
)
(
    input [DATA_WIDTH - 1 : 0] din,
    output [DATA_WIDTH - 1 : 0] dout
);

reg [][] mem;


endmodule;